module UART_rx
(
    clk,
    serialData,
    outputData
);
    